module supersc(	input clk,
						input reset
						
);

endmodule
